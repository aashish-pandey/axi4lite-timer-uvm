class timer_cov extends uvm_component;
    `uvm_component_utils(timer_cov)

    function new(string name="timer_cov", uvm_component parent = null);
        super.new(name, parent);
    endfunction

endclass